module decoder_5to32(in, out);
	input [4:0] in;
	output [31:0] out;
endmodule